LIBRARY IEEE;
USE IEEE.Std_Logic_1164.ALL;

ENTITY MUX_PE IS
	PORT (
		pe_out : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		IR_Out : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		d : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END ENTITY MUX_PE;

ARCHITECTURE arch OF MUX_PE IS
	SIGNAL d_out : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN

	WITH pe_out SELECT
		d_out <= "11111110" WHEN "000",
		"11111101" WHEN "001",
		"11111011" WHEN "010",
		"11110111" WHEN "011",
		"11101111" WHEN "100",
		"11011111" WHEN "101",
		"10111111" WHEN "110",
		"01111111" WHEN OTHERS;
	d <= (IR_Out(15 DOWNTO 8) & d_out) AND IR_Out;
END ARCHITECTURE arch;