LIBRARY IEEE;
USE IEEE.Std_Logic_1164.ALL;

PACKAGE mypkg IS
	TYPE reg_bus IS ARRAY(0 TO 7) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
END PACKAGE mypkg;